// qsys_top.v

// Generated using ACDS version 23.4 66

`timescale 1 ps / 1 ps
module qsys_top (
		input  wire       clk_clk,                          //                       clk.clk
		output wire [3:0] pio_0_external_connection_export  // pio_0_external_connection.export
	);

	wire         clock_in_out_clk_clk;                                           // clock_in:out_clk -> iopll_0:refclk
	wire         iopll_0_outclk0_clk;                                            // iopll_0:outclk_0 -> [intel_niosv_m_0:clk, intel_onchip_memory_0:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:iopll_0_outclk0_clk, pio_0:clk, rst_controller:clk, rst_controller_001:clk, sysid_qsys_0:clock]
	wire         reset_release_0_ninit_done_reset;                               // reset_release_0:ninit_done -> iopll_0:rst
	wire  [31:0] intel_niosv_m_0_data_manager_awaddr;                            // intel_niosv_m_0:data_manager_awaddr -> mm_interconnect_0:intel_niosv_m_0_data_manager_awaddr
	wire   [1:0] intel_niosv_m_0_data_manager_bresp;                             // mm_interconnect_0:intel_niosv_m_0_data_manager_bresp -> intel_niosv_m_0:data_manager_bresp
	wire         intel_niosv_m_0_data_manager_arready;                           // mm_interconnect_0:intel_niosv_m_0_data_manager_arready -> intel_niosv_m_0:data_manager_arready
	wire  [31:0] intel_niosv_m_0_data_manager_rdata;                             // mm_interconnect_0:intel_niosv_m_0_data_manager_rdata -> intel_niosv_m_0:data_manager_rdata
	wire   [3:0] intel_niosv_m_0_data_manager_wstrb;                             // intel_niosv_m_0:data_manager_wstrb -> mm_interconnect_0:intel_niosv_m_0_data_manager_wstrb
	wire         intel_niosv_m_0_data_manager_wready;                            // mm_interconnect_0:intel_niosv_m_0_data_manager_wready -> intel_niosv_m_0:data_manager_wready
	wire         intel_niosv_m_0_data_manager_awready;                           // mm_interconnect_0:intel_niosv_m_0_data_manager_awready -> intel_niosv_m_0:data_manager_awready
	wire         intel_niosv_m_0_data_manager_rready;                            // intel_niosv_m_0:data_manager_rready -> mm_interconnect_0:intel_niosv_m_0_data_manager_rready
	wire         intel_niosv_m_0_data_manager_bready;                            // intel_niosv_m_0:data_manager_bready -> mm_interconnect_0:intel_niosv_m_0_data_manager_bready
	wire         intel_niosv_m_0_data_manager_wvalid;                            // intel_niosv_m_0:data_manager_wvalid -> mm_interconnect_0:intel_niosv_m_0_data_manager_wvalid
	wire  [31:0] intel_niosv_m_0_data_manager_araddr;                            // intel_niosv_m_0:data_manager_araddr -> mm_interconnect_0:intel_niosv_m_0_data_manager_araddr
	wire   [2:0] intel_niosv_m_0_data_manager_arprot;                            // intel_niosv_m_0:data_manager_arprot -> mm_interconnect_0:intel_niosv_m_0_data_manager_arprot
	wire   [1:0] intel_niosv_m_0_data_manager_rresp;                             // mm_interconnect_0:intel_niosv_m_0_data_manager_rresp -> intel_niosv_m_0:data_manager_rresp
	wire   [2:0] intel_niosv_m_0_data_manager_awprot;                            // intel_niosv_m_0:data_manager_awprot -> mm_interconnect_0:intel_niosv_m_0_data_manager_awprot
	wire  [31:0] intel_niosv_m_0_data_manager_wdata;                             // intel_niosv_m_0:data_manager_wdata -> mm_interconnect_0:intel_niosv_m_0_data_manager_wdata
	wire         intel_niosv_m_0_data_manager_arvalid;                           // intel_niosv_m_0:data_manager_arvalid -> mm_interconnect_0:intel_niosv_m_0_data_manager_arvalid
	wire         intel_niosv_m_0_data_manager_bvalid;                            // mm_interconnect_0:intel_niosv_m_0_data_manager_bvalid -> intel_niosv_m_0:data_manager_bvalid
	wire         intel_niosv_m_0_data_manager_awvalid;                           // intel_niosv_m_0:data_manager_awvalid -> mm_interconnect_0:intel_niosv_m_0_data_manager_awvalid
	wire         intel_niosv_m_0_data_manager_rvalid;                            // mm_interconnect_0:intel_niosv_m_0_data_manager_rvalid -> intel_niosv_m_0:data_manager_rvalid
	wire  [31:0] intel_niosv_m_0_instruction_manager_awaddr;                     // intel_niosv_m_0:instruction_manager_awaddr -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_awaddr
	wire   [1:0] intel_niosv_m_0_instruction_manager_bresp;                      // mm_interconnect_0:intel_niosv_m_0_instruction_manager_bresp -> intel_niosv_m_0:instruction_manager_bresp
	wire         intel_niosv_m_0_instruction_manager_arready;                    // mm_interconnect_0:intel_niosv_m_0_instruction_manager_arready -> intel_niosv_m_0:instruction_manager_arready
	wire  [31:0] intel_niosv_m_0_instruction_manager_rdata;                      // mm_interconnect_0:intel_niosv_m_0_instruction_manager_rdata -> intel_niosv_m_0:instruction_manager_rdata
	wire   [3:0] intel_niosv_m_0_instruction_manager_wstrb;                      // intel_niosv_m_0:instruction_manager_wstrb -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_wstrb
	wire         intel_niosv_m_0_instruction_manager_wready;                     // mm_interconnect_0:intel_niosv_m_0_instruction_manager_wready -> intel_niosv_m_0:instruction_manager_wready
	wire         intel_niosv_m_0_instruction_manager_awready;                    // mm_interconnect_0:intel_niosv_m_0_instruction_manager_awready -> intel_niosv_m_0:instruction_manager_awready
	wire         intel_niosv_m_0_instruction_manager_rready;                     // intel_niosv_m_0:instruction_manager_rready -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_rready
	wire         intel_niosv_m_0_instruction_manager_bready;                     // intel_niosv_m_0:instruction_manager_bready -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_bready
	wire         intel_niosv_m_0_instruction_manager_wvalid;                     // intel_niosv_m_0:instruction_manager_wvalid -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_wvalid
	wire  [31:0] intel_niosv_m_0_instruction_manager_araddr;                     // intel_niosv_m_0:instruction_manager_araddr -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_araddr
	wire   [2:0] intel_niosv_m_0_instruction_manager_arprot;                     // intel_niosv_m_0:instruction_manager_arprot -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_arprot
	wire   [1:0] intel_niosv_m_0_instruction_manager_rresp;                      // mm_interconnect_0:intel_niosv_m_0_instruction_manager_rresp -> intel_niosv_m_0:instruction_manager_rresp
	wire   [2:0] intel_niosv_m_0_instruction_manager_awprot;                     // intel_niosv_m_0:instruction_manager_awprot -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_awprot
	wire  [31:0] intel_niosv_m_0_instruction_manager_wdata;                      // intel_niosv_m_0:instruction_manager_wdata -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_wdata
	wire         intel_niosv_m_0_instruction_manager_arvalid;                    // intel_niosv_m_0:instruction_manager_arvalid -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_arvalid
	wire         intel_niosv_m_0_instruction_manager_bvalid;                     // mm_interconnect_0:intel_niosv_m_0_instruction_manager_bvalid -> intel_niosv_m_0:instruction_manager_bvalid
	wire         intel_niosv_m_0_instruction_manager_awvalid;                    // intel_niosv_m_0:instruction_manager_awvalid -> mm_interconnect_0:intel_niosv_m_0_instruction_manager_awvalid
	wire         intel_niosv_m_0_instruction_manager_rvalid;                     // mm_interconnect_0:intel_niosv_m_0_instruction_manager_rvalid -> intel_niosv_m_0:instruction_manager_rvalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;       // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;    // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [1:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_awburst;         // mm_interconnect_0:intel_onchip_memory_0_axi_s1_awburst -> intel_onchip_memory_0:s1_awburst
	wire   [7:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_arlen;           // mm_interconnect_0:intel_onchip_memory_0_axi_s1_arlen -> intel_onchip_memory_0:s1_arlen
	wire   [3:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_wstrb;           // mm_interconnect_0:intel_onchip_memory_0_axi_s1_wstrb -> intel_onchip_memory_0:s1_wstrb
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_wready;          // intel_onchip_memory_0:s1_wready -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_wready
	wire   [1:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_rid;             // intel_onchip_memory_0:s1_rid -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_rid
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_rready;          // mm_interconnect_0:intel_onchip_memory_0_axi_s1_rready -> intel_onchip_memory_0:s1_rready
	wire   [7:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_awlen;           // mm_interconnect_0:intel_onchip_memory_0_axi_s1_awlen -> intel_onchip_memory_0:s1_awlen
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_wvalid;          // mm_interconnect_0:intel_onchip_memory_0_axi_s1_wvalid -> intel_onchip_memory_0:s1_wvalid
	wire  [19:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_araddr;          // mm_interconnect_0:intel_onchip_memory_0_axi_s1_araddr -> intel_onchip_memory_0:s1_araddr
	wire  [31:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_wdata;           // mm_interconnect_0:intel_onchip_memory_0_axi_s1_wdata -> intel_onchip_memory_0:s1_wdata
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_arvalid;         // mm_interconnect_0:intel_onchip_memory_0_axi_s1_arvalid -> intel_onchip_memory_0:s1_arvalid
	wire   [1:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_arid;            // mm_interconnect_0:intel_onchip_memory_0_axi_s1_arid -> intel_onchip_memory_0:s1_arid
	wire  [19:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_awaddr;          // mm_interconnect_0:intel_onchip_memory_0_axi_s1_awaddr -> intel_onchip_memory_0:s1_awaddr
	wire   [1:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_bresp;           // intel_onchip_memory_0:s1_bresp -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_bresp
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_arready;         // intel_onchip_memory_0:s1_arready -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_arready
	wire  [31:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_rdata;           // intel_onchip_memory_0:s1_rdata -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_rdata
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_awready;         // intel_onchip_memory_0:s1_awready -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_awready
	wire   [1:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_arburst;         // mm_interconnect_0:intel_onchip_memory_0_axi_s1_arburst -> intel_onchip_memory_0:s1_arburst
	wire   [2:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_arsize;          // mm_interconnect_0:intel_onchip_memory_0_axi_s1_arsize -> intel_onchip_memory_0:s1_arsize
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_bready;          // mm_interconnect_0:intel_onchip_memory_0_axi_s1_bready -> intel_onchip_memory_0:s1_bready
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_rlast;           // intel_onchip_memory_0:s1_rlast -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_rlast
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_wlast;           // mm_interconnect_0:intel_onchip_memory_0_axi_s1_wlast -> intel_onchip_memory_0:s1_wlast
	wire   [1:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_rresp;           // intel_onchip_memory_0:s1_rresp -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_rresp
	wire   [1:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_awid;            // mm_interconnect_0:intel_onchip_memory_0_axi_s1_awid -> intel_onchip_memory_0:s1_awid
	wire   [1:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_bid;             // intel_onchip_memory_0:s1_bid -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_bid
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_bvalid;          // intel_onchip_memory_0:s1_bvalid -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_bvalid
	wire   [2:0] mm_interconnect_0_intel_onchip_memory_0_axi_s1_awsize;          // mm_interconnect_0:intel_onchip_memory_0_axi_s1_awsize -> intel_onchip_memory_0:s1_awsize
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_awvalid;         // mm_interconnect_0:intel_onchip_memory_0_axi_s1_awvalid -> intel_onchip_memory_0:s1_awvalid
	wire         mm_interconnect_0_intel_onchip_memory_0_axi_s1_rvalid;          // intel_onchip_memory_0:s1_rvalid -> mm_interconnect_0:intel_onchip_memory_0_axi_s1_rvalid
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;          // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;           // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata;            // intel_niosv_m_0:dm_agent_readdata -> mm_interconnect_0:intel_niosv_m_0_dm_agent_readdata
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest;         // intel_niosv_m_0:dm_agent_waitrequest -> mm_interconnect_0:intel_niosv_m_0_dm_agent_waitrequest
	wire  [15:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_address;             // mm_interconnect_0:intel_niosv_m_0_dm_agent_address -> intel_niosv_m_0:dm_agent_address
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_read;                // mm_interconnect_0:intel_niosv_m_0_dm_agent_read -> intel_niosv_m_0:dm_agent_read
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid;       // intel_niosv_m_0:dm_agent_readdatavalid -> mm_interconnect_0:intel_niosv_m_0_dm_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_m_0_dm_agent_write;               // mm_interconnect_0:intel_niosv_m_0_dm_agent_write -> intel_niosv_m_0:dm_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata;           // mm_interconnect_0:intel_niosv_m_0_dm_agent_writedata -> intel_niosv_m_0:dm_agent_writedata
	wire         mm_interconnect_0_pio_0_s1_chipselect;                          // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                            // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                             // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                               // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                           // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata;      // intel_niosv_m_0:timer_sw_agent_readdata -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_readdata
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest;   // intel_niosv_m_0:timer_sw_agent_waitrequest -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_waitrequest
	wire   [5:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address;       // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_address -> intel_niosv_m_0:timer_sw_agent_address
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read;          // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_read -> intel_niosv_m_0:timer_sw_agent_read
	wire   [3:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable;    // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_byteenable -> intel_niosv_m_0:timer_sw_agent_byteenable
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid; // intel_niosv_m_0:timer_sw_agent_readdatavalid -> mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_readdatavalid
	wire         mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write;         // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_write -> intel_niosv_m_0:timer_sw_agent_write
	wire  [31:0] mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata;     // mm_interconnect_0:intel_niosv_m_0_timer_sw_agent_writedata -> intel_niosv_m_0:timer_sw_agent_writedata
	wire         irq_mapper_receiver0_irq;                                       // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [15:0] intel_niosv_m_0_platform_irq_rx_irq;                            // irq_mapper:sender_irq -> intel_niosv_m_0:platform_irq_rx_irq
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [intel_niosv_m_0:reset_reset, intel_onchip_memory_0:reset, irq_mapper:reset, jtag_uart_0:rst_n, pio_0:reset_n, rst_translator:in_reset, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                             // rst_controller:reset_req -> [intel_onchip_memory_0:reset_req, rst_translator:reset_req_in]
	wire         iopll_0_locked_reset;                                           // iopll_0:locked -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> [mm_interconnect_0:intel_niosv_m_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_translator_reset_reset_bridge_in_reset_reset]

	qsys_top_clock_in clock_in (
		.in_clk  (clk_clk),              //   input,  width = 1,  in_clk.clk
		.out_clk (clock_in_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	qsys_top_intel_niosv_m_0 intel_niosv_m_0 (
		.clk                          (iopll_0_outclk0_clk),                                            //   input,   width = 1,                 clk.clk
		.reset_reset                  (rst_controller_reset_out_reset),                                 //   input,   width = 1,               reset.reset
		.platform_irq_rx_irq          (intel_niosv_m_0_platform_irq_rx_irq),                            //   input,  width = 16,     platform_irq_rx.irq
		.instruction_manager_awaddr   (intel_niosv_m_0_instruction_manager_awaddr),                     //  output,  width = 32, instruction_manager.awaddr
		.instruction_manager_awprot   (intel_niosv_m_0_instruction_manager_awprot),                     //  output,   width = 3,                    .awprot
		.instruction_manager_awvalid  (intel_niosv_m_0_instruction_manager_awvalid),                    //  output,   width = 1,                    .awvalid
		.instruction_manager_awready  (intel_niosv_m_0_instruction_manager_awready),                    //   input,   width = 1,                    .awready
		.instruction_manager_wdata    (intel_niosv_m_0_instruction_manager_wdata),                      //  output,  width = 32,                    .wdata
		.instruction_manager_wstrb    (intel_niosv_m_0_instruction_manager_wstrb),                      //  output,   width = 4,                    .wstrb
		.instruction_manager_wvalid   (intel_niosv_m_0_instruction_manager_wvalid),                     //  output,   width = 1,                    .wvalid
		.instruction_manager_wready   (intel_niosv_m_0_instruction_manager_wready),                     //   input,   width = 1,                    .wready
		.instruction_manager_bresp    (intel_niosv_m_0_instruction_manager_bresp),                      //   input,   width = 2,                    .bresp
		.instruction_manager_bvalid   (intel_niosv_m_0_instruction_manager_bvalid),                     //   input,   width = 1,                    .bvalid
		.instruction_manager_bready   (intel_niosv_m_0_instruction_manager_bready),                     //  output,   width = 1,                    .bready
		.instruction_manager_araddr   (intel_niosv_m_0_instruction_manager_araddr),                     //  output,  width = 32,                    .araddr
		.instruction_manager_arprot   (intel_niosv_m_0_instruction_manager_arprot),                     //  output,   width = 3,                    .arprot
		.instruction_manager_arvalid  (intel_niosv_m_0_instruction_manager_arvalid),                    //  output,   width = 1,                    .arvalid
		.instruction_manager_arready  (intel_niosv_m_0_instruction_manager_arready),                    //   input,   width = 1,                    .arready
		.instruction_manager_rdata    (intel_niosv_m_0_instruction_manager_rdata),                      //   input,  width = 32,                    .rdata
		.instruction_manager_rresp    (intel_niosv_m_0_instruction_manager_rresp),                      //   input,   width = 2,                    .rresp
		.instruction_manager_rvalid   (intel_niosv_m_0_instruction_manager_rvalid),                     //   input,   width = 1,                    .rvalid
		.instruction_manager_rready   (intel_niosv_m_0_instruction_manager_rready),                     //  output,   width = 1,                    .rready
		.data_manager_awaddr          (intel_niosv_m_0_data_manager_awaddr),                            //  output,  width = 32,        data_manager.awaddr
		.data_manager_awprot          (intel_niosv_m_0_data_manager_awprot),                            //  output,   width = 3,                    .awprot
		.data_manager_awvalid         (intel_niosv_m_0_data_manager_awvalid),                           //  output,   width = 1,                    .awvalid
		.data_manager_awready         (intel_niosv_m_0_data_manager_awready),                           //   input,   width = 1,                    .awready
		.data_manager_wdata           (intel_niosv_m_0_data_manager_wdata),                             //  output,  width = 32,                    .wdata
		.data_manager_wstrb           (intel_niosv_m_0_data_manager_wstrb),                             //  output,   width = 4,                    .wstrb
		.data_manager_wvalid          (intel_niosv_m_0_data_manager_wvalid),                            //  output,   width = 1,                    .wvalid
		.data_manager_wready          (intel_niosv_m_0_data_manager_wready),                            //   input,   width = 1,                    .wready
		.data_manager_bresp           (intel_niosv_m_0_data_manager_bresp),                             //   input,   width = 2,                    .bresp
		.data_manager_bvalid          (intel_niosv_m_0_data_manager_bvalid),                            //   input,   width = 1,                    .bvalid
		.data_manager_bready          (intel_niosv_m_0_data_manager_bready),                            //  output,   width = 1,                    .bready
		.data_manager_araddr          (intel_niosv_m_0_data_manager_araddr),                            //  output,  width = 32,                    .araddr
		.data_manager_arprot          (intel_niosv_m_0_data_manager_arprot),                            //  output,   width = 3,                    .arprot
		.data_manager_arvalid         (intel_niosv_m_0_data_manager_arvalid),                           //  output,   width = 1,                    .arvalid
		.data_manager_arready         (intel_niosv_m_0_data_manager_arready),                           //   input,   width = 1,                    .arready
		.data_manager_rdata           (intel_niosv_m_0_data_manager_rdata),                             //   input,  width = 32,                    .rdata
		.data_manager_rresp           (intel_niosv_m_0_data_manager_rresp),                             //   input,   width = 2,                    .rresp
		.data_manager_rvalid          (intel_niosv_m_0_data_manager_rvalid),                            //   input,   width = 1,                    .rvalid
		.data_manager_rready          (intel_niosv_m_0_data_manager_rready),                            //  output,   width = 1,                    .rready
		.timer_sw_agent_write         (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write),         //   input,   width = 1,      timer_sw_agent.write
		.timer_sw_agent_writedata     (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata),     //   input,  width = 32,                    .writedata
		.timer_sw_agent_byteenable    (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable),    //   input,   width = 4,                    .byteenable
		.timer_sw_agent_address       (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address),       //   input,   width = 6,                    .address
		.timer_sw_agent_read          (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read),          //   input,   width = 1,                    .read
		.timer_sw_agent_readdata      (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata),      //  output,  width = 32,                    .readdata
		.timer_sw_agent_readdatavalid (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid), //  output,   width = 1,                    .readdatavalid
		.timer_sw_agent_waitrequest   (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest),   //  output,   width = 1,                    .waitrequest
		.dm_agent_write               (mm_interconnect_0_intel_niosv_m_0_dm_agent_write),               //   input,   width = 1,            dm_agent.write
		.dm_agent_writedata           (mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata),           //   input,  width = 32,                    .writedata
		.dm_agent_address             (mm_interconnect_0_intel_niosv_m_0_dm_agent_address),             //   input,  width = 16,                    .address
		.dm_agent_read                (mm_interconnect_0_intel_niosv_m_0_dm_agent_read),                //   input,   width = 1,                    .read
		.dm_agent_readdata            (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata),            //  output,  width = 32,                    .readdata
		.dm_agent_readdatavalid       (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid),       //  output,   width = 1,                    .readdatavalid
		.dm_agent_waitrequest         (mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest)          //  output,   width = 1,                    .waitrequest
	);

	qsys_top_intel_onchip_memory_0 intel_onchip_memory_0 (
		.clk        (iopll_0_outclk0_clk),                                    //   input,   width = 1,   clk1.clk
		.s1_arid    (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arid),    //   input,   width = 2, axi_s1.arid
		.s1_araddr  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_araddr),  //   input,  width = 20,       .araddr
		.s1_arlen   (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arlen),   //   input,   width = 8,       .arlen
		.s1_arsize  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arsize),  //   input,   width = 3,       .arsize
		.s1_arburst (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arburst), //   input,   width = 2,       .arburst
		.s1_arready (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arready), //  output,   width = 1,       .arready
		.s1_arvalid (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arvalid), //   input,   width = 1,       .arvalid
		.s1_awid    (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awid),    //   input,   width = 2,       .awid
		.s1_awaddr  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awaddr),  //   input,  width = 20,       .awaddr
		.s1_awlen   (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awlen),   //   input,   width = 8,       .awlen
		.s1_awsize  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awsize),  //   input,   width = 3,       .awsize
		.s1_awburst (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awburst), //   input,   width = 2,       .awburst
		.s1_awready (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awready), //  output,   width = 1,       .awready
		.s1_awvalid (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awvalid), //   input,   width = 1,       .awvalid
		.s1_rid     (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rid),     //  output,   width = 2,       .rid
		.s1_rdata   (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rdata),   //  output,  width = 32,       .rdata
		.s1_rlast   (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rlast),   //  output,   width = 1,       .rlast
		.s1_rready  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rready),  //   input,   width = 1,       .rready
		.s1_rvalid  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rvalid),  //  output,   width = 1,       .rvalid
		.s1_rresp   (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rresp),   //  output,   width = 2,       .rresp
		.s1_wdata   (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wdata),   //   input,  width = 32,       .wdata
		.s1_wstrb   (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wstrb),   //   input,   width = 4,       .wstrb
		.s1_wlast   (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wlast),   //   input,   width = 1,       .wlast
		.s1_wready  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wready),  //  output,   width = 1,       .wready
		.s1_wvalid  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wvalid),  //   input,   width = 1,       .wvalid
		.s1_bid     (mm_interconnect_0_intel_onchip_memory_0_axi_s1_bid),     //  output,   width = 2,       .bid
		.s1_bresp   (mm_interconnect_0_intel_onchip_memory_0_axi_s1_bresp),   //  output,   width = 2,       .bresp
		.s1_bready  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_bready),  //   input,   width = 1,       .bready
		.s1_bvalid  (mm_interconnect_0_intel_onchip_memory_0_axi_s1_bvalid),  //  output,   width = 1,       .bvalid
		.reset      (rst_controller_reset_out_reset),                         //   input,   width = 1, reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                      //   input,   width = 1,       .reset_req
	);

	qsys_top_iopll_0 iopll_0 (
		.refclk   (clock_in_out_clk_clk),             //   input,  width = 1,  refclk.clk
		.locked   (iopll_0_locked_reset),             //  output,  width = 1,  locked.reset_n
		.rst      (reset_release_0_ninit_done_reset), //   input,  width = 1,   reset.reset
		.outclk_0 (iopll_0_outclk0_clk)               //  output,  width = 1, outclk0.clk
	);

	qsys_top_jtag_uart_0 jtag_uart_0 (
		.clk            (iopll_0_outclk0_clk),                                         //   input,   width = 1,               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //   input,   width = 1,             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //   input,   width = 1, avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //   input,   width = 1,                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //   input,   width = 1,                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //  output,  width = 32,                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //   input,   width = 1,                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //   input,  width = 32,                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //  output,   width = 1,                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //  output,   width = 1,               irq.irq
	);

	qsys_top_pio_0 pio_0 (
		.clk        (iopll_0_outclk0_clk),                   //   input,   width = 1,                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //   input,   width = 1,               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //   input,   width = 2,                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //   input,   width = 1,                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //   input,  width = 32,                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //   input,   width = 1,                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //  output,  width = 32,                    .readdata
		.out_port   (pio_0_external_connection_export)       //  output,   width = 4, external_connection.export
	);

	qsys_top_s10_user_rst_clkgate_0 reset_release_0 (
		.ninit_done (reset_release_0_ninit_done_reset)  //  output,  width = 1, ninit_done.reset
	);

	qsys_top_sysid_qsys_0 sysid_qsys_0 (
		.clock    (iopll_0_outclk0_clk),                                   //   input,   width = 1,           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //   input,   width = 1,         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), //  output,  width = 32, control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //   input,   width = 1,              .address
	);

	qsys_top_altera_mm_interconnect_1920_fimi64y mm_interconnect_0 (
		.jtag_uart_0_avalon_jtag_slave_address                                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),        //  output,   width = 1,                                        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),          //  output,   width = 1,                                                                     .write
		.jtag_uart_0_avalon_jtag_slave_read                                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),           //  output,   width = 1,                                                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata                                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),       //   input,  width = 32,                                                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),      //  output,  width = 32,                                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),    //   input,   width = 1,                                                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),     //  output,   width = 1,                                                                     .chipselect
		.intel_onchip_memory_0_axi_s1_awid                                          (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awid),            //  output,   width = 2,                                         intel_onchip_memory_0_axi_s1.awid
		.intel_onchip_memory_0_axi_s1_awaddr                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awaddr),          //  output,  width = 20,                                                                     .awaddr
		.intel_onchip_memory_0_axi_s1_awlen                                         (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awlen),           //  output,   width = 8,                                                                     .awlen
		.intel_onchip_memory_0_axi_s1_awsize                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awsize),          //  output,   width = 3,                                                                     .awsize
		.intel_onchip_memory_0_axi_s1_awburst                                       (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awburst),         //  output,   width = 2,                                                                     .awburst
		.intel_onchip_memory_0_axi_s1_awvalid                                       (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awvalid),         //  output,   width = 1,                                                                     .awvalid
		.intel_onchip_memory_0_axi_s1_awready                                       (mm_interconnect_0_intel_onchip_memory_0_axi_s1_awready),         //   input,   width = 1,                                                                     .awready
		.intel_onchip_memory_0_axi_s1_wdata                                         (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wdata),           //  output,  width = 32,                                                                     .wdata
		.intel_onchip_memory_0_axi_s1_wstrb                                         (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wstrb),           //  output,   width = 4,                                                                     .wstrb
		.intel_onchip_memory_0_axi_s1_wlast                                         (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wlast),           //  output,   width = 1,                                                                     .wlast
		.intel_onchip_memory_0_axi_s1_wvalid                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wvalid),          //  output,   width = 1,                                                                     .wvalid
		.intel_onchip_memory_0_axi_s1_wready                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_wready),          //   input,   width = 1,                                                                     .wready
		.intel_onchip_memory_0_axi_s1_bid                                           (mm_interconnect_0_intel_onchip_memory_0_axi_s1_bid),             //   input,   width = 2,                                                                     .bid
		.intel_onchip_memory_0_axi_s1_bresp                                         (mm_interconnect_0_intel_onchip_memory_0_axi_s1_bresp),           //   input,   width = 2,                                                                     .bresp
		.intel_onchip_memory_0_axi_s1_bvalid                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_bvalid),          //   input,   width = 1,                                                                     .bvalid
		.intel_onchip_memory_0_axi_s1_bready                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_bready),          //  output,   width = 1,                                                                     .bready
		.intel_onchip_memory_0_axi_s1_arid                                          (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arid),            //  output,   width = 2,                                                                     .arid
		.intel_onchip_memory_0_axi_s1_araddr                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_araddr),          //  output,  width = 20,                                                                     .araddr
		.intel_onchip_memory_0_axi_s1_arlen                                         (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arlen),           //  output,   width = 8,                                                                     .arlen
		.intel_onchip_memory_0_axi_s1_arsize                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arsize),          //  output,   width = 3,                                                                     .arsize
		.intel_onchip_memory_0_axi_s1_arburst                                       (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arburst),         //  output,   width = 2,                                                                     .arburst
		.intel_onchip_memory_0_axi_s1_arvalid                                       (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arvalid),         //  output,   width = 1,                                                                     .arvalid
		.intel_onchip_memory_0_axi_s1_arready                                       (mm_interconnect_0_intel_onchip_memory_0_axi_s1_arready),         //   input,   width = 1,                                                                     .arready
		.intel_onchip_memory_0_axi_s1_rid                                           (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rid),             //   input,   width = 2,                                                                     .rid
		.intel_onchip_memory_0_axi_s1_rdata                                         (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rdata),           //   input,  width = 32,                                                                     .rdata
		.intel_onchip_memory_0_axi_s1_rresp                                         (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rresp),           //   input,   width = 2,                                                                     .rresp
		.intel_onchip_memory_0_axi_s1_rlast                                         (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rlast),           //   input,   width = 1,                                                                     .rlast
		.intel_onchip_memory_0_axi_s1_rvalid                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rvalid),          //   input,   width = 1,                                                                     .rvalid
		.intel_onchip_memory_0_axi_s1_rready                                        (mm_interconnect_0_intel_onchip_memory_0_axi_s1_rready),          //  output,   width = 1,                                                                     .rready
		.sysid_qsys_0_control_slave_address                                         (mm_interconnect_0_sysid_qsys_0_control_slave_address),           //  output,   width = 1,                                           sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                        (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),          //   input,  width = 32,                                                                     .readdata
		.intel_niosv_m_0_dm_agent_address                                           (mm_interconnect_0_intel_niosv_m_0_dm_agent_address),             //  output,  width = 16,                                             intel_niosv_m_0_dm_agent.address
		.intel_niosv_m_0_dm_agent_write                                             (mm_interconnect_0_intel_niosv_m_0_dm_agent_write),               //  output,   width = 1,                                                                     .write
		.intel_niosv_m_0_dm_agent_read                                              (mm_interconnect_0_intel_niosv_m_0_dm_agent_read),                //  output,   width = 1,                                                                     .read
		.intel_niosv_m_0_dm_agent_readdata                                          (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdata),            //   input,  width = 32,                                                                     .readdata
		.intel_niosv_m_0_dm_agent_writedata                                         (mm_interconnect_0_intel_niosv_m_0_dm_agent_writedata),           //  output,  width = 32,                                                                     .writedata
		.intel_niosv_m_0_dm_agent_readdatavalid                                     (mm_interconnect_0_intel_niosv_m_0_dm_agent_readdatavalid),       //   input,   width = 1,                                                                     .readdatavalid
		.intel_niosv_m_0_dm_agent_waitrequest                                       (mm_interconnect_0_intel_niosv_m_0_dm_agent_waitrequest),         //   input,   width = 1,                                                                     .waitrequest
		.pio_0_s1_address                                                           (mm_interconnect_0_pio_0_s1_address),                             //  output,   width = 2,                                                             pio_0_s1.address
		.pio_0_s1_write                                                             (mm_interconnect_0_pio_0_s1_write),                               //  output,   width = 1,                                                                     .write
		.pio_0_s1_readdata                                                          (mm_interconnect_0_pio_0_s1_readdata),                            //   input,  width = 32,                                                                     .readdata
		.pio_0_s1_writedata                                                         (mm_interconnect_0_pio_0_s1_writedata),                           //  output,  width = 32,                                                                     .writedata
		.pio_0_s1_chipselect                                                        (mm_interconnect_0_pio_0_s1_chipselect),                          //  output,   width = 1,                                                                     .chipselect
		.intel_niosv_m_0_timer_sw_agent_address                                     (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_address),       //  output,   width = 6,                                       intel_niosv_m_0_timer_sw_agent.address
		.intel_niosv_m_0_timer_sw_agent_write                                       (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_write),         //  output,   width = 1,                                                                     .write
		.intel_niosv_m_0_timer_sw_agent_read                                        (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_read),          //  output,   width = 1,                                                                     .read
		.intel_niosv_m_0_timer_sw_agent_readdata                                    (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdata),      //   input,  width = 32,                                                                     .readdata
		.intel_niosv_m_0_timer_sw_agent_writedata                                   (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_writedata),     //  output,  width = 32,                                                                     .writedata
		.intel_niosv_m_0_timer_sw_agent_byteenable                                  (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_byteenable),    //  output,   width = 4,                                                                     .byteenable
		.intel_niosv_m_0_timer_sw_agent_readdatavalid                               (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_readdatavalid), //   input,   width = 1,                                                                     .readdatavalid
		.intel_niosv_m_0_timer_sw_agent_waitrequest                                 (mm_interconnect_0_intel_niosv_m_0_timer_sw_agent_waitrequest),   //   input,   width = 1,                                                                     .waitrequest
		.intel_niosv_m_0_data_manager_awaddr                                        (intel_niosv_m_0_data_manager_awaddr),                            //   input,  width = 32,                                         intel_niosv_m_0_data_manager.awaddr
		.intel_niosv_m_0_data_manager_awprot                                        (intel_niosv_m_0_data_manager_awprot),                            //   input,   width = 3,                                                                     .awprot
		.intel_niosv_m_0_data_manager_awvalid                                       (intel_niosv_m_0_data_manager_awvalid),                           //   input,   width = 1,                                                                     .awvalid
		.intel_niosv_m_0_data_manager_awready                                       (intel_niosv_m_0_data_manager_awready),                           //  output,   width = 1,                                                                     .awready
		.intel_niosv_m_0_data_manager_wdata                                         (intel_niosv_m_0_data_manager_wdata),                             //   input,  width = 32,                                                                     .wdata
		.intel_niosv_m_0_data_manager_wstrb                                         (intel_niosv_m_0_data_manager_wstrb),                             //   input,   width = 4,                                                                     .wstrb
		.intel_niosv_m_0_data_manager_wvalid                                        (intel_niosv_m_0_data_manager_wvalid),                            //   input,   width = 1,                                                                     .wvalid
		.intel_niosv_m_0_data_manager_wready                                        (intel_niosv_m_0_data_manager_wready),                            //  output,   width = 1,                                                                     .wready
		.intel_niosv_m_0_data_manager_bresp                                         (intel_niosv_m_0_data_manager_bresp),                             //  output,   width = 2,                                                                     .bresp
		.intel_niosv_m_0_data_manager_bvalid                                        (intel_niosv_m_0_data_manager_bvalid),                            //  output,   width = 1,                                                                     .bvalid
		.intel_niosv_m_0_data_manager_bready                                        (intel_niosv_m_0_data_manager_bready),                            //   input,   width = 1,                                                                     .bready
		.intel_niosv_m_0_data_manager_araddr                                        (intel_niosv_m_0_data_manager_araddr),                            //   input,  width = 32,                                                                     .araddr
		.intel_niosv_m_0_data_manager_arprot                                        (intel_niosv_m_0_data_manager_arprot),                            //   input,   width = 3,                                                                     .arprot
		.intel_niosv_m_0_data_manager_arvalid                                       (intel_niosv_m_0_data_manager_arvalid),                           //   input,   width = 1,                                                                     .arvalid
		.intel_niosv_m_0_data_manager_arready                                       (intel_niosv_m_0_data_manager_arready),                           //  output,   width = 1,                                                                     .arready
		.intel_niosv_m_0_data_manager_rdata                                         (intel_niosv_m_0_data_manager_rdata),                             //  output,  width = 32,                                                                     .rdata
		.intel_niosv_m_0_data_manager_rresp                                         (intel_niosv_m_0_data_manager_rresp),                             //  output,   width = 2,                                                                     .rresp
		.intel_niosv_m_0_data_manager_rvalid                                        (intel_niosv_m_0_data_manager_rvalid),                            //  output,   width = 1,                                                                     .rvalid
		.intel_niosv_m_0_data_manager_rready                                        (intel_niosv_m_0_data_manager_rready),                            //   input,   width = 1,                                                                     .rready
		.intel_niosv_m_0_instruction_manager_awaddr                                 (intel_niosv_m_0_instruction_manager_awaddr),                     //   input,  width = 32,                                  intel_niosv_m_0_instruction_manager.awaddr
		.intel_niosv_m_0_instruction_manager_awprot                                 (intel_niosv_m_0_instruction_manager_awprot),                     //   input,   width = 3,                                                                     .awprot
		.intel_niosv_m_0_instruction_manager_awvalid                                (intel_niosv_m_0_instruction_manager_awvalid),                    //   input,   width = 1,                                                                     .awvalid
		.intel_niosv_m_0_instruction_manager_awready                                (intel_niosv_m_0_instruction_manager_awready),                    //  output,   width = 1,                                                                     .awready
		.intel_niosv_m_0_instruction_manager_wdata                                  (intel_niosv_m_0_instruction_manager_wdata),                      //   input,  width = 32,                                                                     .wdata
		.intel_niosv_m_0_instruction_manager_wstrb                                  (intel_niosv_m_0_instruction_manager_wstrb),                      //   input,   width = 4,                                                                     .wstrb
		.intel_niosv_m_0_instruction_manager_wvalid                                 (intel_niosv_m_0_instruction_manager_wvalid),                     //   input,   width = 1,                                                                     .wvalid
		.intel_niosv_m_0_instruction_manager_wready                                 (intel_niosv_m_0_instruction_manager_wready),                     //  output,   width = 1,                                                                     .wready
		.intel_niosv_m_0_instruction_manager_bresp                                  (intel_niosv_m_0_instruction_manager_bresp),                      //  output,   width = 2,                                                                     .bresp
		.intel_niosv_m_0_instruction_manager_bvalid                                 (intel_niosv_m_0_instruction_manager_bvalid),                     //  output,   width = 1,                                                                     .bvalid
		.intel_niosv_m_0_instruction_manager_bready                                 (intel_niosv_m_0_instruction_manager_bready),                     //   input,   width = 1,                                                                     .bready
		.intel_niosv_m_0_instruction_manager_araddr                                 (intel_niosv_m_0_instruction_manager_araddr),                     //   input,  width = 32,                                                                     .araddr
		.intel_niosv_m_0_instruction_manager_arprot                                 (intel_niosv_m_0_instruction_manager_arprot),                     //   input,   width = 3,                                                                     .arprot
		.intel_niosv_m_0_instruction_manager_arvalid                                (intel_niosv_m_0_instruction_manager_arvalid),                    //   input,   width = 1,                                                                     .arvalid
		.intel_niosv_m_0_instruction_manager_arready                                (intel_niosv_m_0_instruction_manager_arready),                    //  output,   width = 1,                                                                     .arready
		.intel_niosv_m_0_instruction_manager_rdata                                  (intel_niosv_m_0_instruction_manager_rdata),                      //  output,  width = 32,                                                                     .rdata
		.intel_niosv_m_0_instruction_manager_rresp                                  (intel_niosv_m_0_instruction_manager_rresp),                      //  output,   width = 2,                                                                     .rresp
		.intel_niosv_m_0_instruction_manager_rvalid                                 (intel_niosv_m_0_instruction_manager_rvalid),                     //  output,   width = 1,                                                                     .rvalid
		.intel_niosv_m_0_instruction_manager_rready                                 (intel_niosv_m_0_instruction_manager_rready),                     //   input,   width = 1,                                                                     .rready
		.intel_niosv_m_0_reset_reset_bridge_in_reset_reset                          (rst_controller_001_reset_out_reset),                             //   input,   width = 1,                          intel_niosv_m_0_reset_reset_bridge_in_reset.reset
		.jtag_uart_0_avalon_jtag_slave_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                             //   input,   width = 1, jtag_uart_0_avalon_jtag_slave_translator_reset_reset_bridge_in_reset.reset
		.iopll_0_outclk0_clk                                                        (iopll_0_outclk0_clk)                                             //   input,   width = 1,                                                      iopll_0_outclk0.clk
	);

	qsys_top_altera_irq_mapper_2001_ghcid5i irq_mapper (
		.clk           (iopll_0_outclk0_clk),                 //   input,   width = 1,       clk.clk
		.reset         (rst_controller_reset_out_reset),      //   input,   width = 1, clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),            //   input,   width = 1, receiver0.irq
		.sender_irq    (intel_niosv_m_0_platform_irq_rx_irq)  //  output,  width = 16,    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~iopll_0_locked_reset),              //   input,  width = 1, reset_in0.reset
		.clk            (iopll_0_outclk0_clk),                //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~iopll_0_locked_reset),              //   input,  width = 1, reset_in0.reset
		.clk            (iopll_0_outclk0_clk),                //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule

// qsys_top_tb.v

// Generated using ACDS version 23.4 66

`timescale 1 ps / 1 ps
module qsys_top_tb (
	);

	wire    qsys_top_inst_clk_bfm_clk_clk; // qsys_top_inst_clk_bfm:clk -> qsys_top_inst:clk_clk

	qsys_top_inst_clk_bfm_ip qsys_top_inst_clk_bfm (
		.clk (qsys_top_inst_clk_bfm_clk_clk)  //  output,  width = 1, clk.clk
	);

	qsys_top qsys_top_inst (
		.clk_clk                          (qsys_top_inst_clk_bfm_clk_clk), //   input,  width = 1,                       clk.clk
		.pio_0_external_connection_export ()                               //  output,  width = 4, pio_0_external_connection.export
	);

endmodule
